JABALPUR ers or switLOCATED IN MADHYA PRADESH.. CONTAINS MANY LOCATIONS TO VISIT   batch program, specify %%variable instead of
%variable.
Reserved command name
/Loads a program into the upper memory area.

XLOAD   ��  �� ��F2 ��Z�� ^��Y �� ��-[drive:][path]filename [parameters]������pp@  �@���  s�              0 @ 0��   X�  J� ��F2 ��Z�� ���Y X� � 
Enter a choice : rmation
2.Open an existing information
3.Return to main menu
TION     ��  �� ��F2 ��c&��F2���P  ���.� JABALPUR            Jabalpur located in the centre of m.p.                                                                                                                                                                         ��  �� Z� ^��Y �� ��-                                   ���	         �� �`RN:�   r� @ 0��2@�   X�  J� Z� ���Y X� � 
Enter a choice : rmation
2.Open an existing information
3.Return to main menu
TION SYSTEM    ��  �� c&�F2���P  ��Z m,                  n mjkth                                                                                                                                                                                                        ��  �� Z� ^��Y �� ��-                                   ���	         �� �`RN:�   r� @ 0��2@�   X�  J� Z� ���Y X� � 
Enter a choice : rmation
2.Open an existing information
3.Return to main menu
TION SYSTEM    ��  �� c&�F2���P  ��  